`define PARALLEL_ORDER   2
`define PIPELINE_ORDER   1

`define MULT_DATA_WIDTH    32

`define REG_DATA_WIDTH     32
`define REG_ENTRY          32
`define REG_ADDR_WIDTH     $clog2(`REG_ENTRY)
